module led_anode(D,Y); /*��ģ�����ڽ������ 16
������ D ת��Ϊ�˶�����ܵĸ��ε����������
�� Y���Ӷ���� D �ڰ˶�������ϵ���ʾ��
��ν��ʾ������ */
input logic[3:0] D;
output logic[7:0] Y;
always @(D)
begin
case(D)
4'b0000:Y=8'b11000000;
4'b0001:Y=8'b11111001;
4'b0010:Y=8'b10100100;
4'b0011:Y=8'b10110000;
4'b0100:Y=8'b10011001;
4'b0101:Y=8'b10010010;
4'b0110:Y=8'b10000010;
4'b0111:Y=8'b11111000;
4'b1000:Y=8'b10000000;
4'b1001:Y=8'b10010000;
4'b1010:Y=8'b10001000;
4'b1011:Y=8'b10000011;
4'b1100:Y=8'b11000110;
4'b1101:Y=8'b10100001;
4'b1110:Y=8'b10000110;
4'b1111:Y=8'b10001110;
endcase
end
endmodule