`timescale 1ns/1ps
`include"defines.svh"

module openmips_min_sopc(

	input	logic										clk,
	input logic										rst
	
);

  //����ָ��洢��
  InstAddr_t inst_addr;
  Inst_t inst;
  logic rom_ce;
 
 inst_rom inst_rom0(
		.addr(inst_addr),
		.inst(inst),
		.ce(rom_ce)	
	);

 openmips openmips0(
		.clk(clk),
		.rst(rst),
	
		.rom_addr_o(inst_addr),
		.rom_data_i(inst),
		.rom_ce_o(rom_ce)
	
	);
	
	

endmodule